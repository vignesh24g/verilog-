module hello;
	$display(“Hello HDL world”);
end module